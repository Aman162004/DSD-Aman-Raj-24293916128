`timescale 1ns / 1ps

module D_flipflop(
input d, clk,
    output q, qbar
    );
    
 wire sg, rg;

assign #1 sg = ~(clk & d);
assign #1 rg = ~(clk & ~d);
assign #1 q = ~(sg & qbar);
assign #1 qbar = ~(rg & q);

endmodule
