`timescale 1ns / 1ps

module tb_FA(

    );
    
reg A, B, Cin;
wire Sum, Cout;

full_adder uut (
    .A(A),
    .B(B),
    .Cin(Cin),
    .Sum(Sum),
    .Cout(Cout)
);

initial begin
 $dumpfile("dump.vcd");
 $dumpvars(0, tb_FA);

 A=0; B=0; Cin=0; #10;

 A=0; B=0; Cin=1; #10;
    
 A=0; B=1; Cin=0; #10;
 A=0; B=1; Cin=1; #10;
 A=1; B=0; Cin=0; #10;
 A=1; B=0; Cin=1; #10;
 A=1; B=1; Cin=0; #10;
 A=1; B=1; Cin=1; #10;

$finish;
end
endmodule
