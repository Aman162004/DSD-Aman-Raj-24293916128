`timescale 1ns / 1ps


module NOT_gate(
    input a,
    output b
    );
    
assign b = ~a;
    
endmodule
